module main

fn d8p1() int {
    return 0
}

fn d8p2() int {
    return 0
}

fn day8() {
    println('/=== Day 8 ===/')
    println('	- part 1: ${d8p1()}')
    println('	- part 2: ${d8p2()}')
}
