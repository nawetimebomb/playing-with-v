module main

fn d7p1() int {
    return 0
}

fn d7p2() int {
    return 0
}

fn day7() {
    println('/=== Day 7 ===/')
    println('	- part 1: ${d7p1()}')
    println('	- part 2: ${d7p2()}')
}
