module main

fn d14p1() int {
    return 0
}

fn d14p2() int {
    return 0
}

fn day14() {
    println('/=== Day 14 ===/')
    println('	- part 1: ${d14p1()}')
    println('	- part 2: ${d14p2()}')
}
