module main

fn d15p1() int {
    return 0
}

fn d15p2() int {
    return 0
}

fn day15() {
    println('/=== Day 15 ===/')
    println('	- part 1: ${d15p1()}')
    println('	- part 2: ${d15p2()}')
}
