module main

fn part1() int {
    return 0
}

fn part2() int {
    return 0
}

fn main() {
    println('/=== Day 15 ===/')
    println('	- part 1: ${part1()}')
    println('	- part 2: ${part2()}')
}
