module main

fn d5p1() int {
    return 0
}

fn d5p2() int {
    return 0
}

fn day5() {
    println('/=== Day 5 ===/')
    println('	- part 1: ${d5p1()}')
    println('	- part 2: ${d5p2()}')
}
