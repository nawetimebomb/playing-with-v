module main

fn d6p1() int {
    return 0
}

fn d6p2() int {
    return 0
}

fn day6() {
    println('/=== Day 6 ===/')
    println('	- part 1: ${d6p1()}')
    println('	- part 2: ${d6p2()}')
}
