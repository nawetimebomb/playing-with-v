module main

fn d13p1() int {
    return 0
}

fn d13p2() int {
    return 0
}

fn day13() {
    println('/=== Day 13 ===/')
    println('	- part 1: ${d13p1()}')
    println('	- part 2: ${d13p2()}')
}
