module main

fn d10p1() int {
    return 0
}

fn d10p2() int {
    return 0
}

fn day10() {
    println('/=== Day 10 ===/')
    println('	- part 1: ${d10p1()}')
    println('	- part 2: ${d10p2()}')
}
