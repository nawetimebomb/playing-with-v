module main

fn d25p1() int {
    return 0
}

fn d25p2() int {
    return 0
}

fn day25() {
    println('/=== Day 25 ===/')
    println('	- part 1: ${d25p1()}')
    println('	- part 2: ${d25p2()}')
}
