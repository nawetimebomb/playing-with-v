module main

fn d22p1() int {
    return 0
}

fn d22p2() int {
    return 0
}

fn day22() {
    println('/=== Day 22 ===/')
    println('	- part 1: ${d22p1()}')
    println('	- part 2: ${d22p2()}')
}
