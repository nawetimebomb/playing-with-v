module main

fn main() {
	println('Hello, NaweTimebomb')
}
