module main

fn d23p1() int {
    return 0
}

fn d23p2() int {
    return 0
}

fn day23() {
    println('/=== Day 23 ===/')
    println('	- part 1: ${d23p1()}')
    println('	- part 2: ${d23p2()}')
}
