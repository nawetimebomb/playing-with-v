module main

fn d16p1() int {
    return 0
}

fn d16p2() int {
    return 0
}

fn day16() {
    println('/=== Day 16 ===/')
    println('	- part 1: ${d16p1()}')
    println('	- part 2: ${d16p2()}')
}
