module main

fn d4p1() int {
    return 0
}

fn d4p2() int {
    return 0
}

fn day4() {
    println('/=== Day 4 ===/')
    println('	- part 1: ${d4p1()}')
    println('	- part 2: ${d4p2()}')
}
