module main

fn d24p1() int {
    return 0
}

fn d24p2() int {
    return 0
}

fn day24() {
    println('/=== Day 24 ===/')
    println('	- part 1: ${d24p1()}')
    println('	- part 2: ${d24p2()}')
}
