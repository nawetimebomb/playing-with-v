module main

fn d2p1() int {
    return 0
}

fn d2p2() int {
    return 0
}

fn day2() {
    println('/=== Day 2 ===/')
    println('	- part 1: ${d2p1()}')
    println('	- part 2: ${d2p2()}')
}
