module main

fn d3p1() int {
    return 0
}

fn d3p2() int {
    return 0
}

fn day3() {
    println('/=== Day 3 ===/')
    println('	- part 1: ${d3p1()}')
    println('	- part 2: ${d3p2()}')
}
