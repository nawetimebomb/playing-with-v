module main

fn d11p1() int {
    return 0
}

fn d11p2() int {
    return 0
}

fn day11() {
    println('/=== Day 11 ===/')
    println('	- part 1: ${d11p1()}')
    println('	- part 2: ${d11p2()}')
}
