module main

fn d20p1() int {
    return 0
}

fn d20p2() int {
    return 0
}

fn day20() {
    println('/=== Day 20 ===/')
    println('	- part 1: ${d20p1()}')
    println('	- part 2: ${d20p2()}')
}
