module main

fn d19p1() int {
    return 0
}

fn d19p2() int {
    return 0
}

fn day19() {
    println('/=== Day 19 ===/')
    println('	- part 1: ${d19p1()}')
    println('	- part 2: ${d19p2()}')
}
