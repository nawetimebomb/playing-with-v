module main

fn d17p1() int {
    return 0
}

fn d17p2() int {
    return 0
}

fn day17() {
    println('/=== Day 17 ===/')
    println('	- part 1: ${d17p1()}')
    println('	- part 2: ${d17p2()}')
}
