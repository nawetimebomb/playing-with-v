module main

fn d21p1() int {
    return 0
}

fn d21p2() int {
    return 0
}

fn day21() {
    println('/=== Day 21 ===/')
    println('	- part 1: ${d21p1()}')
    println('	- part 2: ${d21p2()}')
}
