module main

fn d9p1() int {
    return 0
}

fn d9p2() int {
    return 0
}

fn day9() {
    println('/=== Day 9 ===/')
    println('	- part 1: ${d9p1()}')
    println('	- part 2: ${d9p2()}')
}
