module main

fn d1p1() int {
    return 0
}

fn d1p2() int {
    return 0
}

fn day1() {
    println('/=== Day 1 ===/')
    println('	- part 1: ${d1p1()}')
    println('	- part 2: ${d1p2()}')
}
