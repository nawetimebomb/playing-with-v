module main

fn d12p1() int {
    return 0
}

fn d12p2() int {
    return 0
}

fn day12() {
    println('/=== Day 12 ===/')
    println('	- part 1: ${d12p1()}')
    println('	- part 2: ${d12p2()}')
}
