module main

fn d18p1() int {
    return 0
}

fn d18p2() int {
    return 0
}

fn day18() {
    println('/=== Day 18 ===/')
    println('	- part 1: ${d18p1()}')
    println('	- part 2: ${d18p2()}')
}
