module main

fn main() {
	day1()
	day2()
}
